Library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
Entity FSM is
	Port(clk,rst :in std_logic;-- Clock and Reset.
		rROM,rRAM,wRAM : out std_logic;--output signals from the FSM.
		Address:out std_logic_vector(1 downto 0));--output Address from the FSM.
End Entity;

Architecture bhv of FSM is
Type FSMType is (S1,S2,S3,S4,S5,S6,S7,S8);--Define an FSM's type.
signal PS : FSMType := S1;--Declare the FSM.
Begin
	Process (clk,rst) is
	Begin
		if rst = '0' Then--If rst is LOW.
			PS <= S1;--reset the FSM.
		Elsif clk'event and clk = '0' Then--On the negative edge.
			--Go the the successor state unconditionally.
			case PS is
				when S1 =>
					PS <= S2;
				when S2 =>
					PS <= S3;
				when S3 =>
					PS <= S4;
				when S4 =>
					PS <= S5;
				when S5 =>
					PS <= S6;
				when S6 =>
					PS <= S7;
				when S7 =>
					PS <= S8;
				when S8 =>
					PS <= S1;
			End Case;
		End if;
	End Process;
	Process (PS)
	Begin
		--Outputs of the FSM depending on the table of the LAB sheet.
		case PS is
			when S1 =>
				Address <= "00";
				rROM <= '1';
				wRAM <= '1';
				rRAM <= '0';
			when S2 =>
				Address <= "01";
				rROM <= '1';
				wRAM <= '1';
				rRAM <= '0';
			when S3 =>
				Address <= "10";
				rROM <= '1';
				wRAM <= '1';
				rRAM <= '0';
			when S4 =>
				Address <= "11";
				rROM <= '1';
				wRAM <= '1';
				rRAM <= '0';
			when S5 =>
				Address <= "00";
				rROM <= '0';
				wRAM <= '0';
				rRAM <= '1';
			when S6 =>
				Address <= "01";
				rROM <= '0';
				wRAM <= '0';
				rRAM <= '1';
			when S7 =>
				Address <= "10";
				rROM <= '0';
				wRAM <= '0';
				rRAM <= '1';
			when S8 =>
				Address <= "11";
				rROM <= '0';
				wRAM <= '0';
				rRAM <= '1';
		End Case;
	End Process;
End;
